----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/10/2025 09:18:46 AM
-- Design Name: 
-- Module Name: edge_detector - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity edge_detector is
    Port ( CLK100MHZ : in STD_LOGIC;
           input : in STD_LOGIC;
           output : out STD_LOGIC);
end edge_detector;

architecture Behavioral of edge_detector is

signal prev_inp : std_logic := '0';
  
begin
        process (CLK100MHZ)
        begin
            if (rising_edge (CLK100MHZ)) then
            
                if (input = '1') then
                    if (prev_inp = '0') then
                        output <= '1';
                    else
                        output <= '0';
                    end if;
                    prev_inp <= '1';
                else    
               
                   prev_inp <= '0';
                
                end if;
                
            end if;
            
                
        end process;

end Behavioral;
